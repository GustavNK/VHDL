library ieee;
use ieee.std_logic_1164.all;

entity Baud_Rate_Generator is
generic(
	
);
	port(
	
);
end;

architecture arch of Baud_Rate_Generator is
begin
	
end;