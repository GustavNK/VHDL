library ieee;
use ieee.std_logic_1164.all;
use work.all;

entity guess_game_test is
port(
	SW	: in std_logic_vector(3 downto 0);
	HEX0	: out std_logic_vector(6 downto 0)
);
end;

architecture guess_game_test_arch of guess_game_test is
begin

end;